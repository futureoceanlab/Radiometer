allan@Allans-MBP-2.local.40852