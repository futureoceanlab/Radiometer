allan@Allans-MBP.local.568